////////////////////////////////////////////////////////////////////////////////
// Sun Aug 17 20:13:33 2025
// Verilog file for RetimeFanout
// naja version: 0.2.5
// Git hash: d4c850b5
////////////////////////////////////////////////////////////////////////////////

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:46.1-92.10" *)
(* top=1 *)
(* hdlname="=RetimeFanout" *)
module RetimeFanout(input clock, input reset, input [15:0] io_in_0, input [15:0] io_in_1,
 output [15:0] io_out);
wire _0000_;
wire _0001_;
wire _0002_;
wire _0003_;
wire _0004_;
wire _0005_;
wire _0006_;
wire _0007_;
wire _0008_;
wire _0009_;
wire _0010_;
wire _0011_;
wire _0012_;
wire _0013_;
wire _0014_;
wire _0015_;
wire _0016_;
wire _0017_;
wire _0018_;
wire _0019_;
wire _0020_;
wire _0021_;
wire _0022_;
wire _0023_;
wire _0024_;
wire _0025_;
wire _0026_;
wire _0027_;
wire _0028_;
wire _0029_;
wire _0030_;
wire _0031_;
wire _0032_;
wire _0033_;
wire _0034_;
wire _0035_;
wire _0036_;
wire _0037_;
wire _0038_;
wire _0039_;
wire _0040_;
wire _0041_;
wire _0042_;
wire _0043_;
wire _0044_;
wire _0045_;
wire _0046_;
wire _0047_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0048_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0049_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0050_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0051_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0052_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0053_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0054_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0055_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0056_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0057_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0058_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0059_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0060_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0061_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0062_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0063_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0064_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0065_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0066_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0067_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0068_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0069_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0070_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0071_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0072_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0073_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0074_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0075_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0076_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0077_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0078_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0079_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0080_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0081_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0082_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0083_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0084_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0085_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0086_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0087_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0088_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0089_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0090_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0091_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0092_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0093_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0094_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0095_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0096_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0097_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0098_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0099_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0100_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0101_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0102_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0103_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0104_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0105_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0106_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0107_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0108_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0109_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0110_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0111_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0112_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0113_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0114_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0115_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0116_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0117_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0118_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0119_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0120_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0121_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0122_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0123_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0124_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0125_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0126_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0127_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0128_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0129_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0130_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0131_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0132_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0133_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0134_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0135_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0136_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0137_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0138_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0139_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0140_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0141_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0142_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0143_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0144_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0145_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0146_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0147_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0148_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0149_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0150_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0151_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0152_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0153_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0154_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0155_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0156_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0157_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0158_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0159_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0160_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0161_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0162_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0163_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0164_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0165_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0166_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0167_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0168_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0169_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0170_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0171_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0172_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0173_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0174_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0175_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0176_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0177_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0178_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0179_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0180_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0181_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0182_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0183_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0184_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0185_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0186_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0187_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0188_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0189_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0190_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0191_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0192_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0193_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0194_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0195_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0196_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0197_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0198_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0199_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0200_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0201_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0202_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0203_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0204_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0205_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0206_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0207_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0208_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0209_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0210_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0211_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0212_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0213_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0214_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0215_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0216_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0217_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0218_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0219_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0220_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0221_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0222_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0223_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0224_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0225_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0226_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0227_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0228_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0229_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0230_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0231_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0232_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0233_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0234_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0235_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0236_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0237_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0238_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0239_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0240_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0241_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0242_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0243_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0244_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0245_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0246_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0247_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0248_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0249_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0250_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0251_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0252_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0253_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0254_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0255_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0256_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0257_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0258_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0259_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0260_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0261_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0262_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0263_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0264_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0265_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0266_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0267_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0268_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0269_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0270_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0271_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0272_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0273_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0274_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0275_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0276_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0277_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0278_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0279_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0280_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0281_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0282_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0283_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0284_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0285_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0286_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0287_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0288_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0289_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0290_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0291_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0292_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0293_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0294_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0295_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0296_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0297_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0298_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0299_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0300_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0301_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0302_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0303_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0304_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0305_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0306_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0307_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0308_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0309_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0310_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0311_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0312_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0313_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0314_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0315_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0316_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0317_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0318_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0319_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0320_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0321_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0322_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0323_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0324_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0325_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0326_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0327_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0328_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0329_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0330_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0331_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0332_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0333_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0334_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0335_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0336_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0337_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0338_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0339_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0340_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0341_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0342_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0343_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0344_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0345_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0346_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0347_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0348_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0349_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0350_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0351_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0352_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0353_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0354_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0355_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0356_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0357_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0358_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0359_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0360_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0361_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0362_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0363_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0364_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0365_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0366_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0367_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0368_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0369_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0370_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0371_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0372_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0373_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0374_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0375_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0376_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0377_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0378_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0379_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0380_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0381_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0382_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0383_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0384_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0385_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0386_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0387_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0388_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0389_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0390_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0391_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0392_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0393_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0394_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0395_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0396_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0397_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0398_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0399_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0400_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0401_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0402_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0403_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0404_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0405_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0406_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0407_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0408_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0409_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0410_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0411_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0412_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0413_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0414_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0415_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0416_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0417_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0418_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0419_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0420_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0421_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0422_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0423_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0424_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0425_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0426_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0427_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0428_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0429_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0430_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0431_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0432_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0433_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0434_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0435_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0436_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0437_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0438_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0439_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0440_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0441_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0442_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0443_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0444_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0445_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0446_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0447_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0448_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0449_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0450_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0451_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0452_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0453_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.26-8.27" *)
wire _0454_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0455_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0456_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0457_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0458_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0459_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0460_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0461_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0462_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0463_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0464_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0465_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0466_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:8.29-8.30" *)
wire _0467_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0468_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0469_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.22-10.24" *)
wire _0470_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:10.26-10.28" *)
wire _0471_;
wire _0472_;
wire _0473_;
wire _0474_;
wire _0475_;
wire _0476_;
wire _0477_;
wire _0478_;
wire _0479_;
wire _0480_;
wire _0481_;
wire _0482_;
wire _0483_;
wire _0484_;
wire _0485_;
wire _0486_;
wire _0487_;
wire _0488_;
wire _0489_;
wire _0490_;
wire _0491_;
wire _0492_;
wire _0493_;
wire _0494_;
wire _0495_;
wire _0496_;
wire _0497_;
wire _0498_;
wire _0499_;
wire _0500_;
wire _0501_;
wire _0502_;
wire _0503_;
wire _0504_;
wire _0505_;
wire _0506_;
wire _0507_;
wire _0508_;
wire _0509_;
wire _0510_;
wire _0511_;
wire _0512_;
wire _0513_;
wire _0514_;
wire _0515_;
wire _0516_;
wire _0517_;
wire _0518_;
wire _0519_;
wire _0520_;
wire _0521_;
wire _0522_;
wire _0523_;
wire _0524_;
wire _0525_;
wire _0526_;
wire _0527_;
wire _0528_;
wire _0529_;
wire _0530_;
wire _0531_;
wire _0532_;
wire _0533_;
wire _0534_;
wire _0535_;
wire _0536_;
wire _0537_;
wire _0538_;
wire _0539_;
wire _0540_;
wire _0541_;
wire _0542_;
wire _0543_;
wire _0544_;
wire _0545_;
wire _0546_;
wire _0547_;
wire _0548_;
wire _0549_;
wire _0550_;
wire _0551_;
wire _0552_;
wire _0553_;
wire _0554_;
wire _0555_;
wire _0556_;
wire _0557_;
wire _0558_;
wire _0559_;
wire _0560_;
wire _0561_;
wire _0562_;
wire _0563_;
wire _0564_;
wire _0565_;
wire _0566_;
wire _0567_;
wire _0568_;
wire _0569_;
wire _0570_;
wire _0571_;
wire _0572_;
wire _0573_;
wire _0574_;
wire _0575_;
wire _0576_;
wire _0577_;
wire _0578_;
wire _0579_;
wire _0580_;
wire _0581_;
wire _0582_;
wire _0583_;
wire _0584_;
wire _0585_;
wire _0586_;
wire _0587_;
wire _0588_;
wire _0589_;
wire _0590_;
wire _0591_;
wire _0592_;
wire _0593_;
wire _0594_;
wire _0595_;
wire _0596_;
wire _0597_;
wire _0598_;
wire _0599_;
wire _0600_;
wire _0601_;
wire _0602_;
wire _0603_;
wire _0604_;
wire _0605_;
wire _0606_;
wire _0607_;
wire _0608_;
wire _0609_;
wire _0610_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0611_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0612_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0613_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0614_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0615_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0616_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0617_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0618_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0619_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0620_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0621_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0622_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0623_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0624_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0625_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0626_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0627_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0628_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0629_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0630_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0631_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0632_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0633_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0634_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0635_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0636_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0637_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0638_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0639_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0640_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0641_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0642_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0643_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0644_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0645_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0646_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0647_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0648_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0649_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0650_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0651_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0652_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0653_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0654_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0655_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0656_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0657_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0658_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0659_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0660_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0661_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0662_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0663_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0664_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0665_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0666_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0667_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0668_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.31-6.32" *)
wire _0669_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0670_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0671_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0672_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0673_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0674_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0675_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0676_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0677_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0678_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0679_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0680_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0681_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0682_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0683_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0684_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0685_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.25-6.26" *)
wire _0686_;
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:6.28-6.29" *)
wire _0687_;

BUFx2_ASAP7_75t_R _0688_ (
  .Y(_0520_),
  .A(io_in_1[0])
);

BUFx2_ASAP7_75t_R _0689_ (
  .Y(_0521_),
  .A(io_in_0[1])
);

AND2x2_ASAP7_75t_R _0690_ (
  .Y(_0289_),
  .A(_0520_),
  .B(_0521_)
);

BUFx2_ASAP7_75t_R _0691_ (
  .Y(_0522_),
  .A(io_in_0[0])
);

BUFx2_ASAP7_75t_R _0692_ (
  .Y(_0523_),
  .A(io_in_1[1])
);

AND2x2_ASAP7_75t_R _0693_ (
  .Y(_0288_),
  .A(_0522_),
  .B(_0523_)
);

BUFx2_ASAP7_75t_R _0694_ (
  .Y(_0524_),
  .A(io_in_0[2])
);

AND2x2_ASAP7_75t_R _0695_ (
  .Y(_0050_),
  .A(io_in_1[0]),
  .B(_0524_)
);

AND2x2_ASAP7_75t_R _0696_ (
  .Y(_0049_),
  .A(_0521_),
  .B(io_in_1[1])
);

BUFx2_ASAP7_75t_R _0697_ (
  .Y(_0525_),
  .A(io_in_1[2])
);

AND2x2_ASAP7_75t_R _0698_ (
  .Y(_0048_),
  .A(_0522_),
  .B(_0525_)
);

BUFx2_ASAP7_75t_R _0699_ (
  .Y(_0526_),
  .A(io_in_0[3])
);

NAND2x1_ASAP7_75t_R _0700_ (
  .Y(_0057_),
  .A(_0520_),
  .B(_0526_)
);

NAND2x1_ASAP7_75t_R _0701_ (
  .Y(_0056_),
  .A(_0523_),
  .B(_0524_)
);

NAND2x1_ASAP7_75t_R _0702_ (
  .Y(_0055_),
  .A(_0521_),
  .B(_0525_)
);

BUFx2_ASAP7_75t_R _0703_ (
  .Y(_0527_),
  .A(io_in_1[3])
);

AND2x2_ASAP7_75t_R _0704_ (
  .Y(_0059_),
  .A(_0522_),
  .B(_0527_)
);

BUFx2_ASAP7_75t_R _0705_ (
  .Y(_0528_),
  .A(io_in_0[4])
);

NAND2x1_ASAP7_75t_R _0706_ (
  .Y(_0066_),
  .A(_0520_),
  .B(_0528_)
);

NAND2x1_ASAP7_75t_R _0707_ (
  .Y(_0065_),
  .A(_0523_),
  .B(_0526_)
);

NAND2x1_ASAP7_75t_R _0708_ (
  .Y(_0064_),
  .A(_0524_),
  .B(_0525_)
);

AND2x2_ASAP7_75t_R _0709_ (
  .Y(_0302_),
  .A(_0521_),
  .B(_0527_)
);

BUFx2_ASAP7_75t_R _0710_ (
  .Y(_0529_),
  .A(io_in_1[4])
);

AND2x2_ASAP7_75t_R _0711_ (
  .Y(_0301_),
  .A(_0522_),
  .B(_0529_)
);

BUFx2_ASAP7_75t_R _0712_ (
  .Y(_0530_),
  .A(io_in_0[5])
);

NAND2x1_ASAP7_75t_R _0713_ (
  .Y(_0072_),
  .A(_0520_),
  .B(_0530_)
);

NAND2x1_ASAP7_75t_R _0714_ (
  .Y(_0071_),
  .A(_0523_),
  .B(_0528_)
);

NAND2x1_ASAP7_75t_R _0715_ (
  .Y(_0070_),
  .A(_0525_),
  .B(_0526_)
);

BUFx2_ASAP7_75t_R _0716_ (
  .Y(_0531_),
  .A(io_in_1[5])
);

NAND2x1_ASAP7_75t_R _0717_ (
  .Y(_0075_),
  .A(_0522_),
  .B(_0531_)
);

BUFx6f_ASAP7_75t_R _0718_ (
  .Y(_0532_),
  .A(io_in_0[6])
);

NAND2x1_ASAP7_75t_R _0719_ (
  .Y(_0085_),
  .A(_0520_),
  .B(_0532_)
);

NAND2x1_ASAP7_75t_R _0720_ (
  .Y(_0084_),
  .A(_0523_),
  .B(_0530_)
);

NAND2x1_ASAP7_75t_R _0721_ (
  .Y(_0083_),
  .A(_0525_),
  .B(_0528_)
);

NAND2x1_ASAP7_75t_R _0722_ (
  .Y(_0089_),
  .A(_0526_),
  .B(_0527_)
);

BUFx6f_ASAP7_75t_R _0723_ (
  .Y(_0533_),
  .A(io_in_1[6])
);

AND2x2_ASAP7_75t_R _0724_ (
  .Y(_0325_),
  .A(_0522_),
  .B(_0533_)
);

BUFx6f_ASAP7_75t_R _0725_ (
  .Y(_0534_),
  .A(io_in_0[8])
);

NAND2x1_ASAP7_75t_R _0726_ (
  .Y(_0096_),
  .A(_0520_),
  .B(_0534_)
);

BUFx6f_ASAP7_75t_R _0727_ (
  .Y(_0535_),
  .A(io_in_0[7])
);

NAND2x1_ASAP7_75t_R _0728_ (
  .Y(_0095_),
  .A(_0523_),
  .B(_0535_)
);

NAND2x1_ASAP7_75t_R _0729_ (
  .Y(_0094_),
  .A(_0525_),
  .B(_0532_)
);

AND2x2_ASAP7_75t_R _0730_ (
  .Y(_0106_),
  .A(io_in_1[1]),
  .B(_0532_)
);

AND2x2_ASAP7_75t_R _0731_ (
  .Y(_0105_),
  .A(io_in_1[2]),
  .B(_0530_)
);

NAND2x1_ASAP7_75t_R _0732_ (
  .Y(_0101_),
  .A(_0527_),
  .B(_0530_)
);

NAND2x1_ASAP7_75t_R _0733_ (
  .Y(_0100_),
  .A(_0528_),
  .B(_0529_)
);

NAND2x1_ASAP7_75t_R _0734_ (
  .Y(_0099_),
  .A(_0526_),
  .B(_0531_)
);

NAND2x1_ASAP7_75t_R _0735_ (
  .Y(_0116_),
  .A(_0524_),
  .B(_0533_)
);

BUFx6f_ASAP7_75t_R _0736_ (
  .Y(_0536_),
  .A(io_in_1[7])
);

NAND2x1_ASAP7_75t_R _0737_ (
  .Y(_0115_),
  .A(_0521_),
  .B(_0536_)
);

BUFx6f_ASAP7_75t_R _0738_ (
  .Y(_0537_),
  .A(io_in_1[8])
);

NAND2x1_ASAP7_75t_R _0739_ (
  .Y(_0114_),
  .A(_0522_),
  .B(_0537_)
);

AND2x2_ASAP7_75t_R _0740_ (
  .Y(_0342_),
  .A(_0521_),
  .B(_0533_)
);

AND2x2_ASAP7_75t_R _0741_ (
  .Y(_0341_),
  .A(_0522_),
  .B(_0536_)
);

BUFx6f_ASAP7_75t_R _0742_ (
  .Y(_0538_),
  .A(io_in_0[9])
);

NAND2x1_ASAP7_75t_R _0743_ (
  .Y(_0133_),
  .A(_0520_),
  .B(_0538_)
);

NAND2x1_ASAP7_75t_R _0744_ (
  .Y(_0134_),
  .A(_0523_),
  .B(_0534_)
);

NAND2x1_ASAP7_75t_R _0745_ (
  .Y(_0132_),
  .A(_0525_),
  .B(_0535_)
);

NAND2x1_ASAP7_75t_R _0746_ (
  .Y(_0139_),
  .A(_0527_),
  .B(_0532_)
);

NAND2x1_ASAP7_75t_R _0747_ (
  .Y(_0138_),
  .A(_0529_),
  .B(_0530_)
);

NAND2x1_ASAP7_75t_R _0748_ (
  .Y(_0137_),
  .A(_0528_),
  .B(_0531_)
);

NAND2x1_ASAP7_75t_R _0749_ (
  .Y(_0145_),
  .A(_0526_),
  .B(_0533_)
);

AND2x2_ASAP7_75t_R _0750_ (
  .Y(_0371_),
  .A(_0522_),
  .B(io_in_1[9])
);

BUFx3_ASAP7_75t_R _0751_ (
  .Y(_0539_),
  .A(io_in_0[10])
);

NAND2x1_ASAP7_75t_R _0752_ (
  .Y(_0151_),
  .A(_0520_),
  .B(_0539_)
);

NAND2x1_ASAP7_75t_R _0753_ (
  .Y(_0150_),
  .A(_0523_),
  .B(_0538_)
);

NAND2x1_ASAP7_75t_R _0754_ (
  .Y(_0152_),
  .A(_0525_),
  .B(_0534_)
);

NAND2x1_ASAP7_75t_R _0755_ (
  .Y(_0157_),
  .A(_0527_),
  .B(_0535_)
);

NAND2x1_ASAP7_75t_R _0756_ (
  .Y(_0155_),
  .A(_0529_),
  .B(_0532_)
);

NAND2x1_ASAP7_75t_R _0757_ (
  .Y(_0156_),
  .A(_0530_),
  .B(_0531_)
);

AND2x2_ASAP7_75t_R _0758_ (
  .Y(_0164_),
  .A(_0526_),
  .B(_0536_)
);

AND2x2_ASAP7_75t_R _0759_ (
  .Y(_0162_),
  .A(_0524_),
  .B(_0537_)
);

AND2x2_ASAP7_75t_R _0760_ (
  .Y(_0390_),
  .A(io_in_0[1]),
  .B(io_in_1[9])
);

AND2x2_ASAP7_75t_R _0761_ (
  .Y(_0389_),
  .A(io_in_0[0]),
  .B(io_in_1[10])
);

INVx1_ASAP7_75t_R _0762_ (
  .Y(_0127_),
  .A(_0470_)
);

NAND2x1_ASAP7_75t_R _0763_ (
  .Y(_0178_),
  .A(_0520_),
  .B(io_in_0[11])
);

NAND2x1_ASAP7_75t_R _0764_ (
  .Y(_0179_),
  .A(_0523_),
  .B(_0539_)
);

NAND2x1_ASAP7_75t_R _0765_ (
  .Y(_0180_),
  .A(_0525_),
  .B(_0538_)
);

NAND2x1_ASAP7_75t_R _0766_ (
  .Y(_0183_),
  .A(_0527_),
  .B(_0534_)
);

NAND2x1_ASAP7_75t_R _0767_ (
  .Y(_0191_),
  .A(_0530_),
  .B(_0533_)
);

NAND2x1_ASAP7_75t_R _0768_ (
  .Y(_0199_),
  .A(_0522_),
  .B(io_in_1[11])
);

NAND2x1_ASAP7_75t_R _0769_ (
  .Y(_0203_),
  .A(_0520_),
  .B(io_in_0[12])
);

AND2x2_ASAP7_75t_R _0770_ (
  .Y(_0208_),
  .A(_0527_),
  .B(_0538_)
);

AND2x2_ASAP7_75t_R _0771_ (
  .Y(_0209_),
  .A(_0529_),
  .B(_0534_)
);

AND2x2_ASAP7_75t_R _0772_ (
  .Y(_0210_),
  .A(_0531_),
  .B(_0535_)
);

AND2x2_ASAP7_75t_R _0773_ (
  .Y(_0213_),
  .A(_0532_),
  .B(_0533_)
);

AND2x2_ASAP7_75t_R _0774_ (
  .Y(_0214_),
  .A(_0530_),
  .B(_0536_)
);

AND2x2_ASAP7_75t_R _0775_ (
  .Y(_0215_),
  .A(_0528_),
  .B(_0537_)
);

AND2x2_ASAP7_75t_R _0776_ (
  .Y(_0220_),
  .A(_0526_),
  .B(io_in_1[9])
);

AND2x2_ASAP7_75t_R _0777_ (
  .Y(_0221_),
  .A(io_in_0[2]),
  .B(io_in_1[10])
);

AND2x2_ASAP7_75t_R _0778_ (
  .Y(_0222_),
  .A(io_in_0[1]),
  .B(io_in_1[11])
);

AND2x2_ASAP7_75t_R _0779_ (
  .Y(_0225_),
  .A(io_in_0[0]),
  .B(io_in_1[12])
);

AND2x2_ASAP7_75t_R _0780_ (
  .Y(_0232_),
  .A(io_in_1[0]),
  .B(io_in_0[13])
);

AND2x2_ASAP7_75t_R _0781_ (
  .Y(_0233_),
  .A(io_in_1[1]),
  .B(io_in_0[12])
);

AND2x2_ASAP7_75t_R _0782_ (
  .Y(_0234_),
  .A(io_in_1[2]),
  .B(io_in_0[11])
);

AND2x2_ASAP7_75t_R _0783_ (
  .Y(_0235_),
  .A(io_in_1[3]),
  .B(_0539_)
);

AND2x2_ASAP7_75t_R _0784_ (
  .Y(_0236_),
  .A(_0529_),
  .B(_0538_)
);

AND2x2_ASAP7_75t_R _0785_ (
  .Y(_0237_),
  .A(_0531_),
  .B(_0534_)
);

AND2x2_ASAP7_75t_R _0786_ (
  .Y(_0240_),
  .A(_0533_),
  .B(_0535_)
);

AND2x2_ASAP7_75t_R _0787_ (
  .Y(_0241_),
  .A(_0532_),
  .B(_0536_)
);

AND2x2_ASAP7_75t_R _0788_ (
  .Y(_0242_),
  .A(_0530_),
  .B(_0537_)
);

AND2x2_ASAP7_75t_R _0789_ (
  .Y(_0246_),
  .A(_0528_),
  .B(io_in_1[9])
);

AND2x2_ASAP7_75t_R _0790_ (
  .Y(_0247_),
  .A(io_in_0[3]),
  .B(io_in_1[10])
);

AND2x2_ASAP7_75t_R _0791_ (
  .Y(_0248_),
  .A(io_in_0[2]),
  .B(io_in_1[11])
);

AND2x2_ASAP7_75t_R _0792_ (
  .Y(_0445_),
  .A(io_in_0[1]),
  .B(io_in_1[12])
);

AND2x2_ASAP7_75t_R _0793_ (
  .Y(_0446_),
  .A(io_in_0[0]),
  .B(io_in_1[13])
);

AND2x2_ASAP7_75t_R _0794_ (
  .Y(_0256_),
  .A(io_in_1[0]),
  .B(io_in_0[14])
);

AND2x2_ASAP7_75t_R _0795_ (
  .Y(_0257_),
  .A(io_in_1[1]),
  .B(io_in_0[13])
);

AND2x2_ASAP7_75t_R _0796_ (
  .Y(_0255_),
  .A(io_in_1[2]),
  .B(io_in_0[12])
);

AND2x2_ASAP7_75t_R _0797_ (
  .Y(_0261_),
  .A(io_in_1[3]),
  .B(io_in_0[11])
);

AND2x2_ASAP7_75t_R _0798_ (
  .Y(_0260_),
  .A(io_in_1[4]),
  .B(_0539_)
);

AND2x2_ASAP7_75t_R _0799_ (
  .Y(_0259_),
  .A(_0531_),
  .B(_0538_)
);

AND2x2_ASAP7_75t_R _0800_ (
  .Y(_0265_),
  .A(_0533_),
  .B(_0534_)
);

AND2x2_ASAP7_75t_R _0801_ (
  .Y(_0266_),
  .A(_0535_),
  .B(_0536_)
);

AND2x2_ASAP7_75t_R _0802_ (
  .Y(_0267_),
  .A(_0532_),
  .B(_0537_)
);

AND2x2_ASAP7_75t_R _0803_ (
  .Y(_0274_),
  .A(_0530_),
  .B(io_in_1[9])
);

AND2x2_ASAP7_75t_R _0804_ (
  .Y(_0275_),
  .A(_0528_),
  .B(io_in_1[10])
);

AND2x2_ASAP7_75t_R _0805_ (
  .Y(_0273_),
  .A(io_in_0[3]),
  .B(io_in_1[11])
);

AND2x2_ASAP7_75t_R _0806_ (
  .Y(_0279_),
  .A(io_in_0[2]),
  .B(io_in_1[12])
);

AND2x2_ASAP7_75t_R _0807_ (
  .Y(_0278_),
  .A(io_in_0[1]),
  .B(io_in_1[13])
);

AND2x2_ASAP7_75t_R _0808_ (
  .Y(_0277_),
  .A(io_in_0[0]),
  .B(io_in_1[14])
);

INVx1_ASAP7_75t_R _0809_ (
  .Y(io_out[9]),
  .A(_0000_)
);

INVx1_ASAP7_75t_R _0810_ (
  .Y(io_out[8]),
  .A(_0001_)
);

INVx1_ASAP7_75t_R _0811_ (
  .Y(io_out[7]),
  .A(_0002_)
);

INVx1_ASAP7_75t_R _0812_ (
  .Y(io_out[6]),
  .A(_0003_)
);

INVx1_ASAP7_75t_R _0813_ (
  .Y(io_out[5]),
  .A(_0004_)
);

INVx1_ASAP7_75t_R _0814_ (
  .Y(io_out[4]),
  .A(_0005_)
);

INVx1_ASAP7_75t_R _0815_ (
  .Y(io_out[3]),
  .A(_0006_)
);

INVx1_ASAP7_75t_R _0816_ (
  .Y(io_out[2]),
  .A(_0007_)
);

INVx1_ASAP7_75t_R _0817_ (
  .Y(io_out[1]),
  .A(_0008_)
);

INVx1_ASAP7_75t_R _0818_ (
  .Y(io_out[15]),
  .A(_0009_)
);

INVx1_ASAP7_75t_R _0819_ (
  .Y(io_out[14]),
  .A(_0010_)
);

INVx1_ASAP7_75t_R _0820_ (
  .Y(io_out[13]),
  .A(_0011_)
);

INVx1_ASAP7_75t_R _0821_ (
  .Y(io_out[12]),
  .A(_0012_)
);

INVx1_ASAP7_75t_R _0822_ (
  .Y(io_out[11]),
  .A(_0013_)
);

INVx1_ASAP7_75t_R _0823_ (
  .Y(io_out[10]),
  .A(_0014_)
);

INVx1_ASAP7_75t_R _0824_ (
  .Y(io_out[0]),
  .A(_0015_)
);

NAND2x1_ASAP7_75t_R _0825_ (
  .Y(_0087_),
  .A(_0521_),
  .B(_0531_)
);

NAND2x1_ASAP7_75t_R _0826_ (
  .Y(_0110_),
  .A(_0524_),
  .B(_0531_)
);

NAND2x1_ASAP7_75t_R _0827_ (
  .Y(_0143_),
  .A(_0521_),
  .B(_0537_)
);

NAND2x1_ASAP7_75t_R _0828_ (
  .Y(_0190_),
  .A(_0526_),
  .B(_0537_)
);

NAND2x1_ASAP7_75t_R _0829_ (
  .Y(_0198_),
  .A(_0521_),
  .B(io_in_1[10])
);

NAND2x1_ASAP7_75t_R _0830_ (
  .Y(_0076_),
  .A(_0521_),
  .B(_0529_)
);

NAND2x1_ASAP7_75t_R _0831_ (
  .Y(_0088_),
  .A(_0524_),
  .B(_0529_)
);

NAND2x1_ASAP7_75t_R _0832_ (
  .Y(_0111_),
  .A(_0526_),
  .B(_0529_)
);

NAND2x1_ASAP7_75t_R _0833_ (
  .Y(_0144_),
  .A(_0524_),
  .B(_0536_)
);

NAND2x1_ASAP7_75t_R _0834_ (
  .Y(_0184_),
  .A(_0529_),
  .B(_0535_)
);

NAND2x1_ASAP7_75t_R _0835_ (
  .Y(_0204_),
  .A(_0523_),
  .B(io_in_0[11])
);

NAND2x1_ASAP7_75t_R _0836_ (
  .Y(_0077_),
  .A(_0524_),
  .B(_0527_)
);

NAND2x1_ASAP7_75t_R _0837_ (
  .Y(_0112_),
  .A(_0527_),
  .B(_0528_)
);

NAND2x1_ASAP7_75t_R _0838_ (
  .Y(_0185_),
  .A(_0531_),
  .B(_0532_)
);

NAND2x1_ASAP7_75t_R _0839_ (
  .Y(_0192_),
  .A(_0528_),
  .B(_0536_)
);

NAND2x1_ASAP7_75t_R _0840_ (
  .Y(_0200_),
  .A(_0524_),
  .B(io_in_1[9])
);

NAND2x1_ASAP7_75t_R _0841_ (
  .Y(_0205_),
  .A(_0525_),
  .B(_0539_)
);

AND2x2_ASAP7_75t_R _0842_ (
  .Y(_0163_),
  .A(io_in_0[4]),
  .B(_0533_)
);

INVx1_ASAP7_75t_R _0843_ (
  .Y(_0175_),
  .A(_0173_)
);

INVx1_ASAP7_75t_R _0844_ (
  .Y(_0398_),
  .A(_0396_)
);

INVx1_ASAP7_75t_R _0845_ (
  .Y(_0434_),
  .A(_0432_)
);

INVx1_ASAP7_75t_R _0846_ (
  .Y(_0397_),
  .A(_0395_)
);

INVx1_ASAP7_75t_R _0847_ (
  .Y(_0455_),
  .A(_0453_)
);

INVx1_ASAP7_75t_R _0848_ (
  .Y(_0284_),
  .A(_0464_)
);

INVx1_ASAP7_75t_R _0849_ (
  .Y(_0467_),
  .A(_0466_)
);

INVx1_ASAP7_75t_R _0850_ (
  .Y(_0336_),
  .A(_0334_)
);

AND2x2_ASAP7_75t_R _0851_ (
  .Y(_0107_),
  .A(io_in_1[0]),
  .B(_0535_)
);

INVx1_ASAP7_75t_R _0852_ (
  .Y(_0351_),
  .A(_0349_)
);

INVx1_ASAP7_75t_R _0853_ (
  .Y(_0379_),
  .A(_0377_)
);

INVx1_ASAP7_75t_R _0854_ (
  .Y(_0176_),
  .A(_0174_)
);

INVx1_ASAP7_75t_R _0855_ (
  .Y(_0378_),
  .A(_0376_)
);

INVx1_ASAP7_75t_R _0856_ (
  .Y(_0416_),
  .A(_0414_)
);

INVx1_ASAP7_75t_R _0857_ (
  .Y(_0417_),
  .A(_0415_)
);

INVx1_ASAP7_75t_R _0858_ (
  .Y(_0433_),
  .A(_0431_)
);

INVx1_ASAP7_75t_R _0859_ (
  .Y(_0454_),
  .A(_0452_)
);

BUFx2_ASAP7_75t_R _0860_ (
  .Y(_0540_),
  .A(reset)
);

INVx1_ASAP7_75t_R _0861_ (
  .Y(_0541_),
  .A(_0540_)
);

AND3x1_ASAP7_75t_R _0862_ (
  .Y(_0472_),
  .A(io_in_1[0]),
  .B(io_in_0[0]),
  .C(_0541_)
);

OA21x2_ASAP7_75t_R _0863_ (
  .Y(_0542_),
  .A1(_0360_),
  .A2(_0470_),
  .B(_0359_)
);

OA21x2_ASAP7_75t_R _0864_ (
  .Y(_0543_),
  .A1(_0381_),
  .A2(_0542_),
  .B(_0380_)
);

XOR2x2_ASAP7_75t_R _0865_ (
  .Y(_0544_),
  .A(_0419_),
  .B(_0543_)
);

AND2x2_ASAP7_75t_R _0866_ (
  .Y(_0473_),
  .A(_0541_),
  .B(_0544_)
);

OA21x2_ASAP7_75t_R _0867_ (
  .Y(_0545_),
  .A1(_0381_),
  .A2(_0130_),
  .B(_0380_)
);

OA21x2_ASAP7_75t_R _0868_ (
  .Y(_0546_),
  .A1(_0419_),
  .A2(_0545_),
  .B(_0418_)
);

XOR2x2_ASAP7_75t_R _0869_ (
  .Y(_0547_),
  .A(_0438_),
  .B(_0546_)
);

AND2x2_ASAP7_75t_R _0870_ (
  .Y(_0474_),
  .A(_0541_),
  .B(_0547_)
);

OA21x2_ASAP7_75t_R _0871_ (
  .Y(_0548_),
  .A1(_0419_),
  .A2(_0543_),
  .B(_0418_)
);

OA21x2_ASAP7_75t_R _0872_ (
  .Y(_0549_),
  .A1(_0438_),
  .A2(_0548_),
  .B(_0437_)
);

XOR2x2_ASAP7_75t_R _0873_ (
  .Y(_0550_),
  .A(_0436_),
  .B(_0549_)
);

AND2x2_ASAP7_75t_R _0874_ (
  .Y(_0475_),
  .A(_0541_),
  .B(_0550_)
);

OA21x2_ASAP7_75t_R _0875_ (
  .Y(_0551_),
  .A1(_0438_),
  .A2(_0546_),
  .B(_0437_)
);

OA21x2_ASAP7_75t_R _0876_ (
  .Y(_0552_),
  .A1(_0436_),
  .A2(_0551_),
  .B(_0435_)
);

XOR2x2_ASAP7_75t_R _0877_ (
  .Y(_0553_),
  .A(_0457_),
  .B(_0552_)
);

AND2x2_ASAP7_75t_R _0878_ (
  .Y(_0476_),
  .A(_0541_),
  .B(_0553_)
);

OR3x1_ASAP7_75t_R _0879_ (
  .Y(_0554_),
  .A(_0436_),
  .B(_0457_),
  .C(_0549_)
);

OA211x2_ASAP7_75t_R _0880_ (
  .Y(_0555_),
  .A1(_0435_),
  .A2(_0457_),
  .B(_0456_),
  .C(_0554_)
);

XOR2x2_ASAP7_75t_R _0881_ (
  .Y(_0556_),
  .A(_0469_),
  .B(_0555_)
);

AND2x2_ASAP7_75t_R _0882_ (
  .Y(_0477_),
  .A(_0541_),
  .B(_0556_)
);

AO21x1_ASAP7_75t_R _0883_ (
  .Y(_0557_),
  .A1(_0457_),
  .A2(_0456_),
  .B(_0469_)
);

AND3x1_ASAP7_75t_R _0884_ (
  .Y(_0558_),
  .A(_0456_),
  .B(_0468_),
  .C(_0552_)
);

AO21x1_ASAP7_75t_R _0885_ (
  .Y(_0559_),
  .A1(_0468_),
  .A2(_0557_),
  .B(_0558_)
);

XOR2x2_ASAP7_75t_R _0886_ (
  .Y(_0560_),
  .A(_0463_),
  .B(_0283_)
);

XNOR2x2_ASAP7_75t_R _0887_ (
  .Y(_0561_),
  .A(_0280_),
  .B(_0285_)
);

XNOR2x2_ASAP7_75t_R _0888_ (
  .Y(_0562_),
  .A(_0560_),
  .B(_0561_)
);

XNOR2x2_ASAP7_75t_R _0889_ (
  .Y(_0563_),
  .A(_0268_),
  .B(_0276_)
);

XNOR2x2_ASAP7_75t_R _0890_ (
  .Y(_0564_),
  .A(_0258_),
  .B(_0262_)
);

XNOR2x2_ASAP7_75t_R _0891_ (
  .Y(_0565_),
  .A(_0563_),
  .B(_0564_)
);

XNOR2x2_ASAP7_75t_R _0892_ (
  .Y(_0566_),
  .A(_0562_),
  .B(_0565_)
);

XOR2x2_ASAP7_75t_R _0893_ (
  .Y(_0567_),
  .A(_0271_),
  .B(_0281_)
);

XNOR2x2_ASAP7_75t_R _0894_ (
  .Y(_0568_),
  .A(_0263_),
  .B(_0269_)
);

XNOR2x2_ASAP7_75t_R _0895_ (
  .Y(_0569_),
  .A(_0567_),
  .B(_0568_)
);

AND2x2_ASAP7_75t_R _0896_ (
  .Y(_0570_),
  .A(io_in_0[2]),
  .B(io_in_1[13])
);

AND2x2_ASAP7_75t_R _0897_ (
  .Y(_0571_),
  .A(io_in_1[3]),
  .B(io_in_0[12])
);

XNOR2x2_ASAP7_75t_R _0898_ (
  .Y(_0572_),
  .A(_0570_),
  .B(_0571_)
);

XNOR2x2_ASAP7_75t_R _0899_ (
  .Y(_0573_),
  .A(_0569_),
  .B(_0572_)
);

XNOR2x2_ASAP7_75t_R _0900_ (
  .Y(_0574_),
  .A(_0566_),
  .B(_0573_)
);

NAND2x1_ASAP7_75t_R _0901_ (
  .Y(_0575_),
  .A(io_in_1[1]),
  .B(io_in_0[14])
);

AND2x2_ASAP7_75t_R _0902_ (
  .Y(_0576_),
  .A(io_in_1[2]),
  .B(io_in_0[13])
);

XNOR2x1_ASAP7_75t_R _0903_ (
  .Y(_0577_),
  .A(_0575_),
  .B(_0576_)
);

AND2x2_ASAP7_75t_R _0904_ (
  .Y(_0578_),
  .A(io_in_1[0]),
  .B(io_in_0[15])
);

AND2x2_ASAP7_75t_R _0905_ (
  .Y(_0579_),
  .A(io_in_1[4]),
  .B(io_in_0[11])
);

XNOR2x1_ASAP7_75t_R _0906_ (
  .Y(_0580_),
  .A(_0578_),
  .B(_0579_)
);

XNOR2x2_ASAP7_75t_R _0907_ (
  .Y(_0581_),
  .A(_0577_),
  .B(_0580_)
);

NAND2x2_ASAP7_75t_R _0908_ (
  .Y(_0582_),
  .A(io_in_0[5]),
  .B(io_in_1[10])
);

AND2x4_ASAP7_75t_R _0909_ (
  .Y(_0583_),
  .A(_0533_),
  .B(_0538_)
);

XNOR2x1_ASAP7_75t_R _0910_ (
  .Y(_0584_),
  .A(_0582_),
  .B(_0583_)
);

AND2x2_ASAP7_75t_R _0911_ (
  .Y(_0585_),
  .A(io_in_0[0]),
  .B(io_in_1[15])
);

AND2x4_ASAP7_75t_R _0912_ (
  .Y(_0586_),
  .A(_0534_),
  .B(_0536_)
);

XNOR2x1_ASAP7_75t_R _0913_ (
  .Y(_0587_),
  .A(_0585_),
  .B(_0586_)
);

XNOR2x1_ASAP7_75t_R _0914_ (
  .Y(_0588_),
  .A(_0584_),
  .B(_0587_)
);

XNOR2x1_ASAP7_75t_R _0915_ (
  .Y(_0589_),
  .A(_0581_),
  .B(_0588_)
);

AND2x2_ASAP7_75t_R _0916_ (
  .Y(_0590_),
  .A(io_in_0[4]),
  .B(io_in_1[11])
);

XOR2x1_ASAP7_75t_R _0917_ (
  .Y(_0591_),
  .A(_0465_),
  .B(_0282_)
);

AND2x2_ASAP7_75t_R _0918_ (
  .Y(_0592_),
  .A(io_in_0[3]),
  .B(io_in_1[12])
);

XNOR2x2_ASAP7_75t_R _0919_ (
  .Y(_0593_),
  .A(_0591_),
  .B(_0592_)
);

XNOR2x1_ASAP7_75t_R _0920_ (
  .Y(_0594_),
  .A(_0590_),
  .B(_0593_)
);

NAND2x1_ASAP7_75t_R _0921_ (
  .Y(_0595_),
  .A(io_in_1[5]),
  .B(_0539_)
);

AND2x4_ASAP7_75t_R _0922_ (
  .Y(_0596_),
  .A(_0535_),
  .B(_0537_)
);

XNOR2x1_ASAP7_75t_R _0923_ (
  .Y(_0597_),
  .A(_0595_),
  .B(_0596_)
);

AND2x2_ASAP7_75t_R _0924_ (
  .Y(_0598_),
  .A(io_in_0[1]),
  .B(io_in_1[14])
);

AND2x4_ASAP7_75t_R _0925_ (
  .Y(_0599_),
  .A(_0532_),
  .B(io_in_1[9])
);

XNOR2x1_ASAP7_75t_R _0926_ (
  .Y(_0600_),
  .A(_0598_),
  .B(_0599_)
);

XNOR2x1_ASAP7_75t_R _0927_ (
  .Y(_0601_),
  .A(_0597_),
  .B(_0600_)
);

XNOR2x1_ASAP7_75t_R _0928_ (
  .Y(_0602_),
  .A(_0594_),
  .B(_0601_)
);

XNOR2x1_ASAP7_75t_R _0929_ (
  .Y(_0603_),
  .A(_0589_),
  .B(_0602_)
);

XNOR2x1_ASAP7_75t_R _0930_ (
  .Y(_0604_),
  .A(_0574_),
  .B(_0603_)
);

XNOR2x1_ASAP7_75t_R _0931_ (
  .Y(_0605_),
  .A(_0559_),
  .B(_0604_)
);

AND2x4_ASAP7_75t_R _0932_ (
  .Y(_0478_),
  .A(_0541_),
  .B(_0605_)
);

BUFx2_ASAP7_75t_R _0933_ (
  .Y(_0606_),
  .A(_0540_)
);

NOR2x1_ASAP7_75t_R _0934_ (
  .Y(_0479_),
  .A(_0606_),
  .B(_0291_)
);

NOR2x1_ASAP7_75t_R _0935_ (
  .Y(_0480_),
  .A(_0606_),
  .B(_0294_)
);

NOR2x1_ASAP7_75t_R _0936_ (
  .Y(_0481_),
  .A(_0606_),
  .B(_0297_)
);

NOR2x1_ASAP7_75t_R _0937_ (
  .Y(_0482_),
  .A(_0606_),
  .B(_0308_)
);

NOR2x1_ASAP7_75t_R _0938_ (
  .Y(_0483_),
  .A(_0606_),
  .B(_0318_)
);

NOR2x1_ASAP7_75t_R _0939_ (
  .Y(_0484_),
  .A(_0606_),
  .B(_0335_)
);

NOR2x1_ASAP7_75t_R _0940_ (
  .Y(_0485_),
  .A(_0606_),
  .B(_0471_)
);

NOR2x1_ASAP7_75t_R _0941_ (
  .Y(_0486_),
  .A(_0606_),
  .B(_0131_)
);

XOR2x2_ASAP7_75t_R _0942_ (
  .Y(_0607_),
  .A(_0381_),
  .B(_0130_)
);

AND2x2_ASAP7_75t_R _0943_ (
  .Y(_0487_),
  .A(_0541_),
  .B(_0607_)
);

BUFx2_ASAP7_75t_R _0944_ (
  .Y(_0608_),
  .A(_0540_)
);

NOR2x1_ASAP7_75t_R _0945_ (
  .Y(_0488_),
  .A(_0047_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0946_ (
  .Y(_0489_),
  .A(_0046_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0947_ (
  .Y(_0490_),
  .A(_0045_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0948_ (
  .Y(_0491_),
  .A(_0044_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0949_ (
  .Y(_0492_),
  .A(_0043_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0950_ (
  .Y(_0493_),
  .A(_0042_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0951_ (
  .Y(_0494_),
  .A(_0041_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0952_ (
  .Y(_0495_),
  .A(_0040_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0953_ (
  .Y(_0496_),
  .A(_0039_),
  .B(_0608_)
);

NOR2x1_ASAP7_75t_R _0954_ (
  .Y(_0497_),
  .A(_0038_),
  .B(_0608_)
);

BUFx2_ASAP7_75t_R _0955_ (
  .Y(_0609_),
  .A(_0540_)
);

NOR2x1_ASAP7_75t_R _0956_ (
  .Y(_0498_),
  .A(_0037_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0957_ (
  .Y(_0499_),
  .A(_0036_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0958_ (
  .Y(_0500_),
  .A(_0035_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0959_ (
  .Y(_0501_),
  .A(_0034_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0960_ (
  .Y(_0502_),
  .A(_0033_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0961_ (
  .Y(_0503_),
  .A(_0032_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0962_ (
  .Y(_0504_),
  .A(_0031_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0963_ (
  .Y(_0505_),
  .A(_0030_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0964_ (
  .Y(_0506_),
  .A(_0029_),
  .B(_0609_)
);

NOR2x1_ASAP7_75t_R _0965_ (
  .Y(_0507_),
  .A(_0028_),
  .B(_0609_)
);

BUFx2_ASAP7_75t_R _0966_ (
  .Y(_0610_),
  .A(_0540_)
);

NOR2x1_ASAP7_75t_R _0967_ (
  .Y(_0508_),
  .A(_0027_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0968_ (
  .Y(_0509_),
  .A(_0026_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0969_ (
  .Y(_0510_),
  .A(_0025_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0970_ (
  .Y(_0511_),
  .A(_0024_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0971_ (
  .Y(_0512_),
  .A(_0023_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0972_ (
  .Y(_0513_),
  .A(_0022_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0973_ (
  .Y(_0514_),
  .A(_0021_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0974_ (
  .Y(_0515_),
  .A(_0020_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0975_ (
  .Y(_0516_),
  .A(_0019_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0976_ (
  .Y(_0517_),
  .A(_0018_),
  .B(_0610_)
);

NOR2x1_ASAP7_75t_R _0977_ (
  .Y(_0518_),
  .A(_0017_),
  .B(_0606_)
);

NOR2x1_ASAP7_75t_R _0978_ (
  .Y(_0519_),
  .A(_0016_),
  .B(_0606_)
);

INVx1_ASAP7_75t_R _0979_ (
  .Y(_0333_),
  .A(_0331_)
);

INVx1_ASAP7_75t_R _0980_ (
  .Y(_0332_),
  .A(_0330_)
);

INVx1_ASAP7_75t_R _0981_ (
  .Y(_0166_),
  .A(_0165_)
);

INVx1_ASAP7_75t_R _0982_ (
  .Y(_0168_),
  .A(_0167_)
);

INVx1_ASAP7_75t_R _0983_ (
  .Y(_0170_),
  .A(_0388_)
);

INVx1_ASAP7_75t_R _0984_ (
  .Y(_0169_),
  .A(_0407_)
);

INVx1_ASAP7_75t_R _0985_ (
  .Y(_0171_),
  .A(_0412_)
);

INVx1_ASAP7_75t_R _0986_ (
  .Y(_0231_),
  .A(_0429_)
);

INVx1_ASAP7_75t_R _0987_ (
  .Y(_0202_),
  .A(_0413_)
);

INVx1_ASAP7_75t_R _0988_ (
  .Y(_0201_),
  .A(_0430_)
);

INVx1_ASAP7_75t_R _0989_ (
  .Y(_0448_),
  .A(_0447_)
);

INVx1_ASAP7_75t_R _0990_ (
  .Y(_0054_),
  .A(_0052_)
);

INVx1_ASAP7_75t_R _0991_ (
  .Y(_0053_),
  .A(_0051_)
);

INVx1_ASAP7_75t_R _0992_ (
  .Y(_0098_),
  .A(_0337_)
);

INVx1_ASAP7_75t_R _0993_ (
  .Y(_0097_),
  .A(_0365_)
);

INVx1_ASAP7_75t_R _0994_ (
  .Y(_0102_),
  .A(_0338_)
);

INVx1_ASAP7_75t_R _0995_ (
  .Y(_0104_),
  .A(_0339_)
);

INVx1_ASAP7_75t_R _0996_ (
  .Y(_0103_),
  .A(_0368_)
);

INVx1_ASAP7_75t_R _0997_ (
  .Y(_0344_),
  .A(_0343_)
);

INVx1_ASAP7_75t_R _0998_ (
  .Y(_0058_),
  .A(_0299_)
);

INVx1_ASAP7_75t_R _0999_ (
  .Y(_0063_),
  .A(_0061_)
);

INVx1_ASAP7_75t_R _1000_ (
  .Y(_0062_),
  .A(_0060_)
);

INVx1_ASAP7_75t_R _1001_ (
  .Y(_0068_),
  .A(_0300_)
);

INVx1_ASAP7_75t_R _1002_ (
  .Y(_0067_),
  .A(_0310_)
);

INVx1_ASAP7_75t_R _1003_ (
  .Y(_0069_),
  .A(_0081_)
);

INVx1_ASAP7_75t_R _1004_ (
  .Y(_0074_),
  .A(_0311_)
);

INVx1_ASAP7_75t_R _1005_ (
  .Y(_0073_),
  .A(_0320_)
);

INVx1_ASAP7_75t_R _1006_ (
  .Y(_0078_),
  .A(_0312_)
);

INVx1_ASAP7_75t_R _1007_ (
  .Y(_0243_),
  .A(_0442_)
);

INVx1_ASAP7_75t_R _1008_ (
  .Y(_0182_),
  .A(_0400_)
);

INVx1_ASAP7_75t_R _1009_ (
  .Y(_0181_),
  .A(_0421_)
);

INVx1_ASAP7_75t_R _1010_ (
  .Y(_0207_),
  .A(_0420_)
);

INVx1_ASAP7_75t_R _1011_ (
  .Y(_0206_),
  .A(_0439_)
);

INVx1_ASAP7_75t_R _1012_ (
  .Y(_0212_),
  .A(_0422_)
);

INVx1_ASAP7_75t_R _1013_ (
  .Y(_0211_),
  .A(_0441_)
);

INVx1_ASAP7_75t_R _1014_ (
  .Y(_0239_),
  .A(_0440_)
);

INVx1_ASAP7_75t_R _1015_ (
  .Y(_0238_),
  .A(_0458_)
);

INVx1_ASAP7_75t_R _1016_ (
  .Y(_0245_),
  .A(_0443_)
);

INVx1_ASAP7_75t_R _1017_ (
  .Y(_0244_),
  .A(_0462_)
);

INVx1_ASAP7_75t_R _1018_ (
  .Y(_0329_),
  .A(_0327_)
);

INVx1_ASAP7_75t_R _1019_ (
  .Y(_0328_),
  .A(_0326_)
);

INVx1_ASAP7_75t_R _1020_ (
  .Y(_0358_),
  .A(_0357_)
);

INVx1_ASAP7_75t_R _1021_ (
  .Y(_0352_),
  .A(_0356_)
);

INVx1_ASAP7_75t_R _1022_ (
  .Y(_0129_),
  .A(_0354_)
);

INVx1_ASAP7_75t_R _1023_ (
  .Y(_0355_),
  .A(_0353_)
);

INVx1_ASAP7_75t_R _1024_ (
  .Y(_0249_),
  .A(_0450_)
);

INVx1_ASAP7_75t_R _1025_ (
  .Y(_0187_),
  .A(_0401_)
);

INVx1_ASAP7_75t_R _1026_ (
  .Y(_0186_),
  .A(_0424_)
);

INVx1_ASAP7_75t_R _1027_ (
  .Y(_0194_),
  .A(_0404_)
);

INVx1_ASAP7_75t_R _1028_ (
  .Y(_0193_),
  .A(_0425_)
);

INVx1_ASAP7_75t_R _1029_ (
  .Y(_0217_),
  .A(_0426_)
);

INVx1_ASAP7_75t_R _1030_ (
  .Y(_0216_),
  .A(_0449_)
);

INVx1_ASAP7_75t_R _1031_ (
  .Y(_0250_),
  .A(_0451_)
);

INVx1_ASAP7_75t_R _1032_ (
  .Y(_0154_),
  .A(_0383_)
);

INVx1_ASAP7_75t_R _1033_ (
  .Y(_0153_),
  .A(_0399_)
);

INVx1_ASAP7_75t_R _1034_ (
  .Y(_0189_),
  .A(_0402_)
);

INVx1_ASAP7_75t_R _1035_ (
  .Y(_0188_),
  .A(_0423_)
);

INVx1_ASAP7_75t_R _1036_ (
  .Y(_0219_),
  .A(_0427_)
);

INVx1_ASAP7_75t_R _1037_ (
  .Y(_0218_),
  .A(_0444_)
);

INVx1_ASAP7_75t_R _1038_ (
  .Y(_0254_),
  .A(_0252_)
);

INVx1_ASAP7_75t_R _1039_ (
  .Y(_0253_),
  .A(_0251_)
);

INVx1_ASAP7_75t_R _1040_ (
  .Y(_0363_),
  .A(_0362_)
);

INVx1_ASAP7_75t_R _1041_ (
  .Y(_0128_),
  .A(_0361_)
);

INVx1_ASAP7_75t_R _1042_ (
  .Y(_0080_),
  .A(_0082_)
);

INVx1_ASAP7_75t_R _1043_ (
  .Y(_0079_),
  .A(_0323_)
);

INVx1_ASAP7_75t_R _1044_ (
  .Y(_0090_),
  .A(_0322_)
);

INVx1_ASAP7_75t_R _1045_ (
  .Y(_0086_),
  .A(_0321_)
);

INVx1_ASAP7_75t_R _1046_ (
  .Y(_0092_),
  .A(_0324_)
);

INVx1_ASAP7_75t_R _1047_ (
  .Y(_0091_),
  .A(_0345_)
);

INVx1_ASAP7_75t_R _1048_ (
  .Y(_0093_),
  .A(_0347_)
);

INVx1_ASAP7_75t_R _1049_ (
  .Y(_0224_),
  .A(_0223_)
);

INVx1_ASAP7_75t_R _1050_ (
  .Y(_0227_),
  .A(_0226_)
);

INVx1_ASAP7_75t_R _1051_ (
  .Y(_0109_),
  .A(_0108_)
);

INVx1_ASAP7_75t_R _1052_ (
  .Y(_0394_),
  .A(_0392_)
);

INVx1_ASAP7_75t_R _1053_ (
  .Y(_0393_),
  .A(_0391_)
);

INVx1_ASAP7_75t_R _1054_ (
  .Y(_0411_),
  .A(_0410_)
);

INVx1_ASAP7_75t_R _1055_ (
  .Y(_0228_),
  .A(_0409_)
);

INVx1_ASAP7_75t_R _1056_ (
  .Y(_0230_),
  .A(_0229_)
);

INVx1_ASAP7_75t_R _1057_ (
  .Y(_0264_),
  .A(_0459_)
);

INVx1_ASAP7_75t_R _1058_ (
  .Y(_0270_),
  .A(_0460_)
);

INVx1_ASAP7_75t_R _1059_ (
  .Y(_0272_),
  .A(_0461_)
);

INVx1_ASAP7_75t_R _1060_ (
  .Y(_0292_),
  .A(_0290_)
);

INVx1_ASAP7_75t_R _1061_ (
  .Y(_0295_),
  .A(_0293_)
);

INVx1_ASAP7_75t_R _1062_ (
  .Y(_0298_),
  .A(_0296_)
);

INVx1_ASAP7_75t_R _1063_ (
  .Y(_0309_),
  .A(_0307_)
);

INVx1_ASAP7_75t_R _1064_ (
  .Y(_0319_),
  .A(_0317_)
);

INVx1_ASAP7_75t_R _1065_ (
  .Y(_0287_),
  .A(_0286_)
);

INVx1_ASAP7_75t_R _1066_ (
  .Y(_0126_),
  .A(_0346_)
);

INVx1_ASAP7_75t_R _1067_ (
  .Y(_0123_),
  .A(_0124_)
);

INVx1_ASAP7_75t_R _1068_ (
  .Y(_0113_),
  .A(_0120_)
);

INVx1_ASAP7_75t_R _1069_ (
  .Y(_0117_),
  .A(_0119_)
);

INVx1_ASAP7_75t_R _1070_ (
  .Y(_0118_),
  .A(_0340_)
);

INVx1_ASAP7_75t_R _1071_ (
  .Y(_0122_),
  .A(_0125_)
);

INVx1_ASAP7_75t_R _1072_ (
  .Y(_0121_),
  .A(_0369_)
);

INVx1_ASAP7_75t_R _1073_ (
  .Y(_0136_),
  .A(_0364_)
);

INVx1_ASAP7_75t_R _1074_ (
  .Y(_0135_),
  .A(_0382_)
);

INVx1_ASAP7_75t_R _1075_ (
  .Y(_0159_),
  .A(_0384_)
);

INVx1_ASAP7_75t_R _1076_ (
  .Y(_0158_),
  .A(_0405_)
);

INVx1_ASAP7_75t_R _1077_ (
  .Y(_0161_),
  .A(_0385_)
);

INVx1_ASAP7_75t_R _1078_ (
  .Y(_0160_),
  .A(_0403_)
);

INVx1_ASAP7_75t_R _1079_ (
  .Y(_0195_),
  .A(_0406_)
);

INVx1_ASAP7_75t_R _1080_ (
  .Y(_0197_),
  .A(_0408_)
);

INVx1_ASAP7_75t_R _1081_ (
  .Y(_0196_),
  .A(_0428_)
);

INVx1_ASAP7_75t_R _1082_ (
  .Y(_0172_),
  .A(_0177_)
);

INVx1_ASAP7_75t_R _1083_ (
  .Y(_0140_),
  .A(_0366_)
);

INVx1_ASAP7_75t_R _1084_ (
  .Y(_0306_),
  .A(_0304_)
);

INVx1_ASAP7_75t_R _1085_ (
  .Y(_0305_),
  .A(_0303_)
);

INVx1_ASAP7_75t_R _1086_ (
  .Y(_0316_),
  .A(_0314_)
);

INVx1_ASAP7_75t_R _1087_ (
  .Y(_0315_),
  .A(_0313_)
);

INVx1_ASAP7_75t_R _1088_ (
  .Y(_0375_),
  .A(_0373_)
);

INVx1_ASAP7_75t_R _1089_ (
  .Y(_0374_),
  .A(_0372_)
);

INVx1_ASAP7_75t_R _1090_ (
  .Y(_0142_),
  .A(_0367_)
);

INVx1_ASAP7_75t_R _1091_ (
  .Y(_0141_),
  .A(_0386_)
);

INVx1_ASAP7_75t_R _1092_ (
  .Y(_0350_),
  .A(_0348_)
);

INVx1_ASAP7_75t_R _1093_ (
  .Y(_0147_),
  .A(_0146_)
);

INVx1_ASAP7_75t_R _1094_ (
  .Y(_0149_),
  .A(_0370_)
);

INVx1_ASAP7_75t_R _1095_ (
  .Y(_0148_),
  .A(_0387_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1096_ (
  .CON(_0051_),
  .SN(_0052_),
  .A(_0048_),
  .B(_0049_),
  .CI(_0050_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1097_ (
  .CON(_0299_),
  .SN(_0611_),
  .A(_0055_),
  .B(_0056_),
  .CI(_0057_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1098_ (
  .CON(_0060_),
  .SN(_0061_),
  .A(_0059_),
  .B(_0053_),
  .CI(_0611_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1099_ (
  .CON(_0310_),
  .SN(_0300_),
  .A(_0064_),
  .B(_0065_),
  .CI(_0066_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1100_ (
  .CON(_0081_),
  .SN(_0670_),
  .A(_0612_),
  .B(_0058_),
  .CI(_0068_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1101_ (
  .CON(_0320_),
  .SN(_0311_),
  .A(_0070_),
  .B(_0071_),
  .CI(_0072_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1102_ (
  .CON(_0672_),
  .SN(_0312_),
  .A(_0075_),
  .B(_0076_),
  .CI(_0077_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1103_ (
  .CON(_0323_),
  .SN(_0082_),
  .A(_0078_),
  .B(_0067_),
  .CI(_0074_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1104_ (
  .CON(_0674_),
  .SN(_0671_),
  .A(_0069_),
  .B(_0080_),
  .CI(_0613_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1105_ (
  .CON(_0619_),
  .SN(_0321_),
  .A(_0083_),
  .B(_0084_),
  .CI(_0085_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1106_ (
  .CON(_0675_),
  .SN(_0322_),
  .A(_0087_),
  .B(_0088_),
  .CI(_0089_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1107_ (
  .CON(_0345_),
  .SN(_0324_),
  .A(_0090_),
  .B(_0073_),
  .CI(_0086_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1108_ (
  .CON(_0347_),
  .SN(_0673_),
  .A(_0614_),
  .B(_0079_),
  .CI(_0092_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1109_ (
  .CON(_0365_),
  .SN(_0337_),
  .A(_0094_),
  .B(_0095_),
  .CI(_0096_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1110_ (
  .CON(_0624_),
  .SN(_0338_),
  .A(_0099_),
  .B(_0100_),
  .CI(_0101_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1111_ (
  .CON(_0368_),
  .SN(_0339_),
  .A(_0102_),
  .B(_0615_),
  .CI(_0098_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1112_ (
  .CON(_0615_),
  .SN(_0108_),
  .A(_0105_),
  .B(_0106_),
  .CI(_0107_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1113_ (
  .CON(_0120_),
  .SN(_0618_),
  .A(_0110_),
  .B(_0111_),
  .CI(_0112_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1114_ (
  .CON(_0626_),
  .SN(_0119_),
  .A(_0114_),
  .B(_0115_),
  .CI(_0116_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1115_ (
  .CON(_0679_),
  .SN(_0340_),
  .A(_0616_),
  .B(_0117_),
  .CI(_0113_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1116_ (
  .CON(_0369_),
  .SN(_0125_),
  .A(_0118_),
  .B(_0617_),
  .CI(_0104_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1117_ (
  .CON(_0617_),
  .SN(_0622_),
  .A(_0618_),
  .B(_0619_),
  .CI(_0109_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1118_ (
  .CON(_0680_),
  .SN(_0677_),
  .A(_0620_),
  .B(_0123_),
  .CI(_0122_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1119_ (
  .CON(_0124_),
  .SN(_0346_),
  .A(_0621_),
  .B(_0091_),
  .CI(_0622_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1120_ (
  .CON(_0676_),
  .SN(_0678_),
  .A(_0623_),
  .B(_0126_),
  .CI(_0093_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1121_ (
  .CON(_0130_),
  .SN(_0131_),
  .A(_0127_),
  .B(_0128_),
  .CI(_0129_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1122_ (
  .CON(_0382_),
  .SN(_0364_),
  .A(_0132_),
  .B(_0133_),
  .CI(_0134_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1123_ (
  .CON(_0630_),
  .SN(_0366_),
  .A(_0137_),
  .B(_0138_),
  .CI(_0139_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1124_ (
  .CON(_0386_),
  .SN(_0367_),
  .A(_0136_),
  .B(_0140_),
  .CI(_0097_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1125_ (
  .CON(_0629_),
  .SN(_0625_),
  .A(_0143_),
  .B(_0144_),
  .CI(_0145_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1126_ (
  .CON(_0146_),
  .SN(_0627_),
  .A(_0624_),
  .B(_0625_),
  .CI(_0626_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1127_ (
  .CON(_0387_),
  .SN(_0370_),
  .A(_0627_),
  .B(_0142_),
  .CI(_0103_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1128_ (
  .CON(_0633_),
  .SN(_0681_),
  .A(_0121_),
  .B(_0628_),
  .CI(_0149_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1129_ (
  .CON(_0399_),
  .SN(_0383_),
  .A(_0150_),
  .B(_0151_),
  .CI(_0152_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1130_ (
  .CON(_0405_),
  .SN(_0384_),
  .A(_0155_),
  .B(_0156_),
  .CI(_0157_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1131_ (
  .CON(_0403_),
  .SN(_0385_),
  .A(_0159_),
  .B(_0135_),
  .CI(_0154_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1132_ (
  .CON(_0635_),
  .SN(_0165_),
  .A(_0162_),
  .B(_0163_),
  .CI(_0164_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1133_ (
  .CON(_0167_),
  .SN(_0631_),
  .A(_0166_),
  .B(_0629_),
  .CI(_0630_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1134_ (
  .CON(_0407_),
  .SN(_0388_),
  .A(_0161_),
  .B(_0141_),
  .CI(_0631_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1135_ (
  .CON(_0412_),
  .SN(_0634_),
  .A(_0632_),
  .B(_0148_),
  .CI(_0170_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1136_ (
  .CON(_0173_),
  .SN(_0174_),
  .A(_0633_),
  .B(_0172_),
  .CI(_0634_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1137_ (
  .CON(_0421_),
  .SN(_0400_),
  .A(_0178_),
  .B(_0179_),
  .CI(_0180_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1138_ (
  .CON(_0424_),
  .SN(_0401_),
  .A(_0183_),
  .B(_0184_),
  .CI(_0185_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1139_ (
  .CON(_0423_),
  .SN(_0402_),
  .A(_0153_),
  .B(_0182_),
  .CI(_0187_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1140_ (
  .CON(_0425_),
  .SN(_0404_),
  .A(_0190_),
  .B(_0191_),
  .CI(_0192_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1141_ (
  .CON(_0641_),
  .SN(_0406_),
  .A(_0194_),
  .B(_0635_),
  .CI(_0158_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1142_ (
  .CON(_0428_),
  .SN(_0408_),
  .A(_0195_),
  .B(_0189_),
  .CI(_0160_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1143_ (
  .CON(_0640_),
  .SN(_0682_),
  .A(_0198_),
  .B(_0199_),
  .CI(_0200_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1144_ (
  .CON(_0430_),
  .SN(_0413_),
  .A(_0169_),
  .B(_0197_),
  .CI(_0636_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1145_ (
  .CON(_0685_),
  .SN(_0683_),
  .A(_0637_),
  .B(_0171_),
  .CI(_0202_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1146_ (
  .CON(_0439_),
  .SN(_0420_),
  .A(_0203_),
  .B(_0204_),
  .CI(_0205_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1147_ (
  .CON(_0646_),
  .SN(_0638_),
  .A(_0208_),
  .B(_0209_),
  .CI(_0210_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1148_ (
  .CON(_0441_),
  .SN(_0422_),
  .A(_0207_),
  .B(_0181_),
  .CI(_0638_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1149_ (
  .CON(_0648_),
  .SN(_0639_),
  .A(_0213_),
  .B(_0214_),
  .CI(_0215_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1150_ (
  .CON(_0449_),
  .SN(_0426_),
  .A(_0186_),
  .B(_0639_),
  .CI(_0193_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1151_ (
  .CON(_0444_),
  .SN(_0427_),
  .A(_0212_),
  .B(_0188_),
  .CI(_0217_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1152_ (
  .CON(_0650_),
  .SN(_0223_),
  .A(_0220_),
  .B(_0221_),
  .CI(_0222_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1153_ (
  .CON(_0652_),
  .SN(_0226_),
  .A(_0224_),
  .B(_0640_),
  .CI(_0225_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1154_ (
  .CON(_0229_),
  .SN(_0642_),
  .A(_0641_),
  .B(_0227_),
  .CI(_0228_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1155_ (
  .CON(_0654_),
  .SN(_0429_),
  .A(_0219_),
  .B(_0196_),
  .CI(_0642_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1156_ (
  .CON(_0686_),
  .SN(_0684_),
  .A(_0231_),
  .B(_0201_),
  .CI(_0643_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1157_ (
  .CON(_0655_),
  .SN(_0644_),
  .A(_0232_),
  .B(_0233_),
  .CI(_0234_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1158_ (
  .CON(_0658_),
  .SN(_0645_),
  .A(_0235_),
  .B(_0236_),
  .CI(_0237_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1159_ (
  .CON(_0458_),
  .SN(_0440_),
  .A(_0644_),
  .B(_0206_),
  .CI(_0645_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1160_ (
  .CON(_0660_),
  .SN(_0647_),
  .A(_0240_),
  .B(_0241_),
  .CI(_0242_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1161_ (
  .CON(_0666_),
  .SN(_0442_),
  .A(_0646_),
  .B(_0647_),
  .CI(_0648_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1162_ (
  .CON(_0462_),
  .SN(_0443_),
  .A(_0239_),
  .B(_0211_),
  .CI(_0243_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1163_ (
  .CON(_0663_),
  .SN(_0649_),
  .A(_0246_),
  .B(_0247_),
  .CI(_0248_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1164_ (
  .CON(_0664_),
  .SN(_0450_),
  .A(_0649_),
  .B(_0650_),
  .CI(_0651_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1165_ (
  .CON(_0687_),
  .SN(_0451_),
  .A(_0216_),
  .B(_0249_),
  .CI(_0652_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1166_ (
  .CON(_0669_),
  .SN(_0653_),
  .A(_0245_),
  .B(_0218_),
  .CI(_0250_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1167_ (
  .CON(_0251_),
  .SN(_0252_),
  .A(_0653_),
  .B(_0230_),
  .CI(_0654_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1168_ (
  .CON(_0258_),
  .SN(_0656_),
  .A(_0255_),
  .B(_0256_),
  .CI(_0257_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1169_ (
  .CON(_0262_),
  .SN(_0657_),
  .A(_0259_),
  .B(_0260_),
  .CI(_0261_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1170_ (
  .CON(_0263_),
  .SN(_0459_),
  .A(_0655_),
  .B(_0656_),
  .CI(_0657_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1171_ (
  .CON(_0268_),
  .SN(_0659_),
  .A(_0265_),
  .B(_0266_),
  .CI(_0267_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1172_ (
  .CON(_0269_),
  .SN(_0460_),
  .A(_0658_),
  .B(_0659_),
  .CI(_0660_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1173_ (
  .CON(_0271_),
  .SN(_0461_),
  .A(_0238_),
  .B(_0264_),
  .CI(_0270_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1174_ (
  .CON(_0276_),
  .SN(_0662_),
  .A(_0273_),
  .B(_0274_),
  .CI(_0275_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1175_ (
  .CON(_0280_),
  .SN(_0661_),
  .A(_0277_),
  .B(_0278_),
  .CI(_0279_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1176_ (
  .CON(_0281_),
  .SN(_0665_),
  .A(_0661_),
  .B(_0662_),
  .CI(_0663_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1177_ (
  .CON(_0282_),
  .SN(_0667_),
  .A(_0664_),
  .B(_0665_),
  .CI(_0666_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1178_ (
  .CON(_0283_),
  .SN(_0668_),
  .A(_0272_),
  .B(_0244_),
  .CI(_0667_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:44.26-46.12" *)
FAx1_ASAP7_75t_R _1179_ (
  .CON(_0285_),
  .SN(_0286_),
  .A(_0668_),
  .B(_0284_),
  .CI(_0669_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1180_ (
  .CON(_0290_),
  .SN(_0291_),
  .A(_0288_),
  .B(_0289_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1181_ (
  .CON(_0293_),
  .SN(_0294_),
  .A(_0292_),
  .B(_0054_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1182_ (
  .CON(_0296_),
  .SN(_0297_),
  .A(_0295_),
  .B(_0063_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1183_ (
  .CON(_0613_),
  .SN(_0612_),
  .A(_0301_),
  .B(_0302_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1184_ (
  .CON(_0303_),
  .SN(_0304_),
  .A(_0062_),
  .B(_0670_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1185_ (
  .CON(_0307_),
  .SN(_0308_),
  .A(_0298_),
  .B(_0306_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1186_ (
  .CON(_0313_),
  .SN(_0314_),
  .A(_0305_),
  .B(_0671_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1187_ (
  .CON(_0317_),
  .SN(_0318_),
  .A(_0309_),
  .B(_0316_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1188_ (
  .CON(_0623_),
  .SN(_0614_),
  .A(_0325_),
  .B(_0672_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1189_ (
  .CON(_0326_),
  .SN(_0327_),
  .A(_0673_),
  .B(_0674_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1190_ (
  .CON(_0330_),
  .SN(_0331_),
  .A(_0315_),
  .B(_0329_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1191_ (
  .CON(_0334_),
  .SN(_0335_),
  .A(_0319_),
  .B(_0333_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1192_ (
  .CON(_0616_),
  .SN(_0343_),
  .A(_0341_),
  .B(_0342_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1193_ (
  .CON(_0620_),
  .SN(_0621_),
  .A(_0344_),
  .B(_0675_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1194_ (
  .CON(_0348_),
  .SN(_0349_),
  .A(_0676_),
  .B(_0677_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1195_ (
  .CON(_0353_),
  .SN(_0354_),
  .A(_0352_),
  .B(_0351_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1196_ (
  .CON(_0356_),
  .SN(_0357_),
  .A(_0328_),
  .B(_0678_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1197_ (
  .CON(_0359_),
  .SN(_0360_),
  .A(_0128_),
  .B(_0129_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1198_ (
  .CON(_0361_),
  .SN(_0362_),
  .A(_0358_),
  .B(_0332_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1199_ (
  .CON(_0177_),
  .SN(_0628_),
  .A(_0371_),
  .B(_0679_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1200_ (
  .CON(_0372_),
  .SN(_0373_),
  .A(_0680_),
  .B(_0681_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1201_ (
  .CON(_0376_),
  .SN(_0377_),
  .A(_0350_),
  .B(_0375_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1202_ (
  .CON(_0380_),
  .SN(_0381_),
  .A(_0355_),
  .B(_0379_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1203_ (
  .CON(_0391_),
  .SN(_0392_),
  .A(_0389_),
  .B(_0390_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1204_ (
  .CON(_0637_),
  .SN(_0632_),
  .A(_0394_),
  .B(_0147_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1205_ (
  .CON(_0395_),
  .SN(_0396_),
  .A(_0374_),
  .B(_0176_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1206_ (
  .CON(_0409_),
  .SN(_0410_),
  .A(_0393_),
  .B(_0682_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1207_ (
  .CON(_0643_),
  .SN(_0636_),
  .A(_0411_),
  .B(_0168_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1208_ (
  .CON(_0414_),
  .SN(_0415_),
  .A(_0175_),
  .B(_0683_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1209_ (
  .CON(_0418_),
  .SN(_0419_),
  .A(_0398_),
  .B(_0378_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1210_ (
  .CON(_0431_),
  .SN(_0432_),
  .A(_0684_),
  .B(_0685_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1211_ (
  .CON(_0435_),
  .SN(_0436_),
  .A(_0434_),
  .B(_0416_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1212_ (
  .CON(_0437_),
  .SN(_0438_),
  .A(_0397_),
  .B(_0417_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1213_ (
  .CON(_0447_),
  .SN(_0651_),
  .A(_0445_),
  .B(_0446_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1214_ (
  .CON(_0452_),
  .SN(_0453_),
  .A(_0686_),
  .B(_0254_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1215_ (
  .CON(_0456_),
  .SN(_0457_),
  .A(_0455_),
  .B(_0433_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1216_ (
  .CON(_0463_),
  .SN(_0464_),
  .A(_0448_),
  .B(_0687_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1217_ (
  .CON(_0465_),
  .SN(_0466_),
  .A(_0287_),
  .B(_0253_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1218_ (
  .CON(_0468_),
  .SN(_0469_),
  .A(_0467_),
  .B(_0454_)
);

(* module_not_derived=32'b00000000000000000000000000000001 *)
(* src="=external/bazel-orfs++orfs_repositories+docker_orfs/OpenROAD-flow-scripts/flow/platforms/asap7/yoSys/cells_adders_R.v:20.29-24.14" *)
HAxp5_ASAP7_75t_R _1219_ (
  .CON(_0470_),
  .SN(_0471_),
  .A(_0336_),
  .B(_0363_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[0]$_SDFF_PP0_  (
  .QN(_0047_),
  .CLK(clock),
  .D(_0472_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[10]$_SDFF_PP0_  (
  .QN(_0046_),
  .CLK(clock),
  .D(_0473_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[11]$_SDFF_PP0_  (
  .QN(_0045_),
  .CLK(clock),
  .D(_0474_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[12]$_SDFF_PP0_  (
  .QN(_0044_),
  .CLK(clock),
  .D(_0475_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[13]$_SDFF_PP0_  (
  .QN(_0043_),
  .CLK(clock),
  .D(_0476_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[14]$_SDFF_PP0_  (
  .QN(_0042_),
  .CLK(clock),
  .D(_0477_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[15]$_SDFF_PP0_  (
  .QN(_0041_),
  .CLK(clock),
  .D(_0478_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[1]$_SDFF_PP0_  (
  .QN(_0040_),
  .CLK(clock),
  .D(_0479_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[2]$_SDFF_PP0_  (
  .QN(_0039_),
  .CLK(clock),
  .D(_0480_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[3]$_SDFF_PP0_  (
  .QN(_0038_),
  .CLK(clock),
  .D(_0481_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[4]$_SDFF_PP0_  (
  .QN(_0037_),
  .CLK(clock),
  .D(_0482_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[5]$_SDFF_PP0_  (
  .QN(_0036_),
  .CLK(clock),
  .D(_0483_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[6]$_SDFF_PP0_  (
  .QN(_0035_),
  .CLK(clock),
  .D(_0484_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[7]$_SDFF_PP0_  (
  .QN(_0034_),
  .CLK(clock),
  .D(_0485_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[8]$_SDFF_PP0_  (
  .QN(_0033_),
  .CLK(clock),
  .D(_0486_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r[9]$_SDFF_PP0_  (
  .QN(_0032_),
  .CLK(clock),
  .D(_0487_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[0]$_SDFF_PP0_  (
  .QN(_0031_),
  .CLK(clock),
  .D(_0488_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[10]$_SDFF_PP0_  (
  .QN(_0030_),
  .CLK(clock),
  .D(_0489_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[11]$_SDFF_PP0_  (
  .QN(_0029_),
  .CLK(clock),
  .D(_0490_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[12]$_SDFF_PP0_  (
  .QN(_0028_),
  .CLK(clock),
  .D(_0491_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[13]$_SDFF_PP0_  (
  .QN(_0027_),
  .CLK(clock),
  .D(_0492_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[14]$_SDFF_PP0_  (
  .QN(_0026_),
  .CLK(clock),
  .D(_0493_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[15]$_SDFF_PP0_  (
  .QN(_0025_),
  .CLK(clock),
  .D(_0494_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[1]$_SDFF_PP0_  (
  .QN(_0024_),
  .CLK(clock),
  .D(_0495_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[2]$_SDFF_PP0_  (
  .QN(_0023_),
  .CLK(clock),
  .D(_0496_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[3]$_SDFF_PP0_  (
  .QN(_0022_),
  .CLK(clock),
  .D(_0497_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[4]$_SDFF_PP0_  (
  .QN(_0021_),
  .CLK(clock),
  .D(_0498_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[5]$_SDFF_PP0_  (
  .QN(_0020_),
  .CLK(clock),
  .D(_0499_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[6]$_SDFF_PP0_  (
  .QN(_0019_),
  .CLK(clock),
  .D(_0500_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[7]$_SDFF_PP0_  (
  .QN(_0018_),
  .CLK(clock),
  .D(_0501_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[8]$_SDFF_PP0_  (
  .QN(_0017_),
  .CLK(clock),
  .D(_0502_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_1[9]$_SDFF_PP0_  (
  .QN(_0016_),
  .CLK(clock),
  .D(_0503_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[0]$_SDFF_PP0_  (
  .QN(_0015_),
  .CLK(clock),
  .D(_0504_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[10]$_SDFF_PP0_  (
  .QN(_0014_),
  .CLK(clock),
  .D(_0505_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[11]$_SDFF_PP0_  (
  .QN(_0013_),
  .CLK(clock),
  .D(_0506_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[12]$_SDFF_PP0_  (
  .QN(_0012_),
  .CLK(clock),
  .D(_0507_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[13]$_SDFF_PP0_  (
  .QN(_0011_),
  .CLK(clock),
  .D(_0508_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[14]$_SDFF_PP0_  (
  .QN(_0010_),
  .CLK(clock),
  .D(_0509_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[15]$_SDFF_PP0_  (
  .QN(_0009_),
  .CLK(clock),
  .D(_0510_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[1]$_SDFF_PP0_  (
  .QN(_0008_),
  .CLK(clock),
  .D(_0511_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[2]$_SDFF_PP0_  (
  .QN(_0007_),
  .CLK(clock),
  .D(_0512_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[3]$_SDFF_PP0_  (
  .QN(_0006_),
  .CLK(clock),
  .D(_0513_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[4]$_SDFF_PP0_  (
  .QN(_0005_),
  .CLK(clock),
  .D(_0514_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[5]$_SDFF_PP0_  (
  .QN(_0004_),
  .CLK(clock),
  .D(_0515_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[6]$_SDFF_PP0_  (
  .QN(_0003_),
  .CLK(clock),
  .D(_0516_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[7]$_SDFF_PP0_  (
  .QN(_0002_),
  .CLK(clock),
  .D(_0517_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[8]$_SDFF_PP0_  (
  .QN(_0001_),
  .CLK(clock),
  .D(_0518_)
);

(* src="=bazel-out/k8-fastbuild/bin/RetimeFanout.sv:57.3-68.6" *)
DFFHQNx1_ASAP7_75t_R \io_out_r_2[9]$_SDFF_PP0_  (
  .QN(_0000_),
  .CLK(clock),
  .D(_0519_)
);
endmodule //RetimeFanout
